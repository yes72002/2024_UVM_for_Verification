`include "uvm_macros.svh"
import uvm_pkg::*;

class spi_config extends uvm_object;  // configuration of env
  `uvm_object_utils(spi_config)

  function new(string name = "spi_config");
    super.new(name);
  endfunction

  uvm_active_passive_enum is_active = UVM_ACTIVE;
endclass

typedef enum bit [1:0] {
  readd  = 0,
  writed = 1,
  rstdut = 2
} oper_mode;

class transaction extends uvm_sequence_item;
  randc logic [7:0] addr;
  rand logic [7:0] din;
  logic [7:0] dout;
  rand oper_mode op;
  logic rst;
  rand logic miso;
  logic cs;
  logic done;
  logic err;
  logic ready;
  logic mosi;

  constraint addr_c {addr <= 10;}

  `uvm_object_utils_begin(transaction)
    `uvm_field_int(addr, UVM_ALL_ON)
    `uvm_field_int(din, UVM_ALL_ON)
    `uvm_field_int(dout, UVM_ALL_ON)
    `uvm_field_int(ready, UVM_ALL_ON)
    `uvm_field_int(rst, UVM_ALL_ON)
    `uvm_field_int(done, UVM_ALL_ON)
    `uvm_field_int(miso, UVM_ALL_ON)
    `uvm_field_int(mosi, UVM_ALL_ON)
    `uvm_field_int(cs, UVM_ALL_ON)
    `uvm_field_int(err, UVM_ALL_ON)
    `uvm_field_enum(oper_mode, op, UVM_DEFAULT)
  `uvm_object_utils_end

  function new(string name = "transaction");
    super.new(name);
  endfunction
endclass : transaction

// write seq
class write_data extends uvm_sequence #(transaction);
  `uvm_object_utils(write_data)

  transaction tr;

  function new(string name = "write_data");
    super.new(name);
  endfunction

  virtual task body();
    repeat (15) begin
      tr = transaction::type_id::create("tr");
      tr.addr_c.constraint_mode(1);
      start_item(tr);
      assert (tr.randomize);
      tr.op = writed;
      finish_item(tr);
    end
  endtask
endclass

class read_data extends uvm_sequence #(transaction);
  `uvm_object_utils(read_data)

  transaction tr;

  function new(string name = "read_data");
    super.new(name);
  endfunction

  virtual task body();
    repeat (15) begin
      tr = transaction::type_id::create("tr");
      tr.addr_c.constraint_mode(1);
      start_item(tr);
      assert (tr.randomize);
      tr.op = readd;
      finish_item(tr);
    end
  endtask
endclass

class reset_dut extends uvm_sequence #(transaction);
  `uvm_object_utils(reset_dut)

  transaction tr;

  function new(string name = "reset_dut");
    super.new(name);
  endfunction

  virtual task body();
    repeat (15) begin
      tr = transaction::type_id::create("tr");
      tr.addr_c.constraint_mode(1);
      start_item(tr);
      assert (tr.randomize);
      tr.op = rstdut;
      finish_item(tr);
    end
  endtask
endclass

class writeb_readb extends uvm_sequence #(transaction);
  `uvm_object_utils(writeb_readb)

  transaction tr;

  function new(string name = "writeb_readb");
    super.new(name);
  endfunction

  virtual task body();
    repeat (10) begin
      tr = transaction::type_id::create("tr");
      tr.addr_c.constraint_mode(1);
      start_item(tr);
      assert (tr.randomize);
      tr.op = writed;
      finish_item(tr);
    end

    repeat (10) begin
      tr = transaction::type_id::create("tr");
      tr.addr_c.constraint_mode(1);
      start_item(tr);
      assert (tr.randomize);
      tr.op = readd;
      finish_item(tr);
    end
  endtask
endclass

class driver extends uvm_driver #(transaction);
  `uvm_component_utils(driver)

  // now working with the driver is a bit tricky
  // We need to get assistance of an interface and hence we add an interface.
  virtual spi_i vif;
  // the trasaction where we will be storing the data that we receive from a sequencer
  transaction tr;
  // data, which is a variable that is capable of holding 16 bits of data.
  logic [15:0] data;  // <- din , addr ->
  logic [7:0] datard;

  function new(input string path = "drv", uvm_component parent = null);
    super.new(path, parent);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    tr = transaction::type_id::create("tr");

    if (!uvm_config_db#(virtual spi_i)::get(this, "", "vif", vif))  // uvm_test_top.env.agent.drv.aif
      `uvm_error("drv", "Unable to access Interface");
  endfunction

  // reset task
  task reset_dut();
    begin
      vif.rst  <= 1'b1;  // active high reset
      vif.miso <= 1'b0;
      vif.cs   <= 1'b1;
      `uvm_info("DRV", "System Reset", UVM_MEDIUM);
      @(posedge vif.clk);
    end
  endtask

  // write
  task write_d();
    // start of transaction, remove the reset
    vif.rst  <= 1'b0;
    vif.cs   <= 1'b0;
    vif.miso <= 1'b0;
    data = {tr.din, tr.addr};
    `uvm_info("DRV", $sformatf("DATA WRITE addr : %0d din : %0d", tr.addr, tr.din), UVM_MEDIUM);
    @(posedge vif.clk);
    vif.miso <= 1'b1;  // write operation
    @(posedge vif.clk);
    for (int i = 0; i < 16; i++) begin
      vif.miso <= data[i];
      @(posedge vif.clk);
    end

    @(posedge vif.op_done);
  endtask

  // read operation
  task read_d();
    // start of transaction, remove the reset
    vif.rst  <= 1'b0;
    vif.cs   <= 1'b0;
    vif.miso <= 1'b0;

    // prepare the data to send
    data = {8'h00, tr.addr};

    @(posedge vif.clk);
    vif.miso <= 1'b0;  // read operation

    // send address
    @(posedge vif.clk);
    for (int i = 0; i < 8; i++) begin
      vif.miso <= data[i];
      // send data in each clock edge
      @(posedge vif.clk);
    end

    // wait for data ready
    @(posedge vif.ready);

    // sample the output data
    for (int i = 0; i < 8; i++) begin
      @(posedge vif.clk);
      datard[i] = vif.mosi;
    end

    // wait for our operation done
    `uvm_info("DRV", $sformatf("DATA READ addr : %0d dout : %0d", tr.addr, datard), UVM_MEDIUM);
    @(posedge vif.op_done);
  endtask

  virtual task run_phase(uvm_phase phase);
    forever begin
      seq_item_port.get_next_item(tr);
      if (tr.op == rstdut) begin
        reset_dut();
      end else if (tr.op == writed) begin
        write_d();
      end else if (tr.op == readd) begin
        read_d();
      end
      seq_item_port.item_done();
    end
  endtask
endclass

class mon extends uvm_monitor;
  `uvm_component_utils(mon)

  uvm_analysis_port #(transaction) send;
  transaction tr;
  virtual spi_i vif;
  logic [15:0] din;
  logic [7:0] dout;

  function new(input string inst = "mon", uvm_component parent = null);
    super.new(inst, parent);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    tr   = transaction::type_id::create("tr");
    send = new("send", this);
    if (!uvm_config_db#(virtual spi_i)::get(this, "", "vif", vif))  //uvm_test_top.env.agent.drv.aif
      `uvm_error("MON", "Unable to access Interface");
  endfunction

  virtual task run_phase(uvm_phase phase);
    forever begin
      @(posedge vif.clk);
      if (vif.rst) begin
        tr.op = rstdut;
        `uvm_info("MON", "SYSTEM RESET DETECTED", UVM_NONE);
        send.write(tr);
      end else begin
        // we will wait for two clock tick (edge) and then check whether chip select (CS)
        // is low and miso is high.
        @(posedge vif.clk);
        if (vif.miso && !vif.cs) begin // write operation
          tr.op = writed;
          @(posedge vif.clk);

          for (int i = 0; i < 16; i++) begin
            din[i] <= vif.miso;
            @(posedge vif.clk);
          end
          // this data will be helpful for a scorebaord to perfrom a comparisoin.
          tr.addr = din[7:0];
          tr.din  = din[15:8];

          @(posedge vif.op_done);
          `uvm_info("MON", $sformatf("DATA WRITE addr:%0d data:%0d", din[7:0], din[15:8]),
                    UVM_NONE);
          send.write(tr);
        end else if (!vif.miso && !vif.cs) begin // read operation
          tr.op = readd;
          @(posedge vif.clk);

          for (int i = 0; i < 8; i++) begin
            din[i] <= vif.miso;
            @(posedge vif.clk);
          end
          tr.addr = din[7:0];

          @(posedge vif.ready);

          for (int i = 0; i < 8; i++) begin
            @(posedge vif.clk);
            dout[i] = vif.mosi;
          end
          @(posedge vif.op_done);
          tr.dout = dout;
          `uvm_info("MON", $sformatf("DATA READ addr:%0d data:%0d ", tr.addr, tr.dout), UVM_NONE);
          send.write(tr);
        end
      end
    end
  endtask
endclass

class sco extends uvm_scoreboard;
  `uvm_component_utils(sco)

  uvm_analysis_imp#(transaction,sco) recv;
  bit [31:0] arr[32] = '{default:0};
  bit [31:0] addr    = 0;
  bit [31:0] data_rd = 0;

  function new(input string inst = "sco", uvm_component parent = null);
    super.new(inst, parent);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    recv = new("recv", this);
  endfunction

  virtual function void write(transaction tr);
    if (tr.op == rstdut) begin
      `uvm_info("SCO", "SYSTEM RESET DETECTED", UVM_NONE);
    end else if (tr.op == writed) begin
      arr[tr.addr] = tr.din;
      `uvm_info("SCO", $sformatf("DATA WRITE OP  addr:%0d, wdata:%0d arr_wr:%0d", tr.addr, tr.din, arr[tr.addr]), UVM_NONE);
    end else if (tr.op == readd) begin
      data_rd = arr[tr.addr];
      if (data_rd == tr.dout)
        `uvm_info(
          "SCO",
          $sformatf("DATA MATCHED : addr:%0d, rdata:%0d", tr.addr, tr.dout),
          UVM_NONE
        )
      else
        `uvm_info(
          "SCO", $sformatf(
          "TEST FAILED : addr:%0d, rdata:%0d data_rd_arr:%0d", tr.addr, tr.dout, data_rd),
          UVM_NONE
        )
    end

    $display("----------------------------------------------------------------");
  endfunction
endclass

class agent extends uvm_agent;
  `uvm_component_utils(agent)

  spi_config cfg;

  function new(input string inst = "agent", uvm_component parent = null);
    super.new(inst, parent);
  endfunction

  driver d;
  uvm_sequencer #(transaction) seqr;
  mon m;

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    cfg = spi_config::type_id::create("cfg");
    m   = mon::type_id::create("m", this);

    if (cfg.is_active == UVM_ACTIVE) begin
      d = driver::type_id::create("d", this);
      seqr = uvm_sequencer#(transaction)::type_id::create("seqr", this);
    end
  endfunction

  virtual function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);
    if (cfg.is_active == UVM_ACTIVE) begin
      d.seq_item_port.connect(seqr.seq_item_export);
    end
  endfunction
endclass

class env extends uvm_env;
  `uvm_component_utils(env)

  function new(input string inst = "env", uvm_component c);
    super.new(inst, c);
  endfunction

  agent a;
  sco   s;

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    a = agent::type_id::create("a", this);
    s = sco::type_id::create("s", this);
  endfunction

  virtual function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);
    a.m.send.connect(s.recv);
  endfunction
endclass

class test extends uvm_test;
  `uvm_component_utils(test)

  function new(input string inst = "test", uvm_component c);
    super.new(inst, c);
  endfunction

  env e;
  write_data wdata;
  read_data rdata;
  writeb_readb wrrdb;
  reset_dut rstdut;

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    e      = env::type_id::create("env", this);
    wdata  = write_data::type_id::create("wdata");
    rdata  = read_data::type_id::create("rdata");
    wrrdb  = writeb_readb::type_id::create("wrrdb");
    rstdut = reset_dut::type_id::create("rstdut");
  endfunction

  virtual task run_phase(uvm_phase phase);
    phase.raise_objection(this);
    wrrdb.start(e.a.seqr);
    phase.drop_objection(this);
  endtask
endclass

module tb;
  spi_i vif ();
  spi_mem dut (
      .clk(vif.clk),
      .rst(vif.rst),
      .cs(vif.cs),
      .miso(vif.miso),
      .ready(vif.ready),
      .mosi(vif.mosi),
      .op_done(vif.op_done)
  );

  initial begin
    vif.clk <= 0;
  end

  always #10 vif.clk <= ~vif.clk;

  initial begin
    uvm_config_db#(virtual spi_i)::set(null, "*", "vif", vif);
    run_test("test");
  end

  initial begin
    $dumpfile("dump.vcd");
    $dumpvars;
  end
endmodule


// # KERNEL: ASDB file was created in location /home/runner/dataset.asdb
// # KERNEL: UVM_INFO @ 0: reporter [RNTST] Running test test...
// # KERNEL: UVM_INFO /home/runner/testbench.sv(190) @ 0: uvm_test_top.env.a.d [DRV] DATA WRITE addr : 4 din : 115
// # KERNEL: UVM_INFO /home/runner/testbench.sv(291) @ 370: uvm_test_top.env.a.m [MON] DATA WRITE addr:4 data:115
// # KERNEL: UVM_INFO /home/runner/testbench.sv(341) @ 370: uvm_test_top.env.s [SCO] DATA WRITE OP  addr:4, wdata:115 arr_wr:115
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/runner/testbench.sv(190) @ 370: uvm_test_top.env.a.d [DRV] DATA WRITE addr : 8 din : 132
// # KERNEL: UVM_INFO /home/runner/testbench.sv(291) @ 750: uvm_test_top.env.a.m [MON] DATA WRITE addr:8 data:132
// # KERNEL: UVM_INFO /home/runner/testbench.sv(341) @ 750: uvm_test_top.env.s [SCO] DATA WRITE OP  addr:8, wdata:132 arr_wr:132
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/runner/testbench.sv(190) @ 750: uvm_test_top.env.a.d [DRV] DATA WRITE addr : 6 din : 166
// # KERNEL: UVM_INFO /home/runner/testbench.sv(291) @ 1130: uvm_test_top.env.a.m [MON] DATA WRITE addr:6 data:166
// # KERNEL: UVM_INFO /home/runner/testbench.sv(341) @ 1130: uvm_test_top.env.s [SCO] DATA WRITE OP  addr:6, wdata:166 arr_wr:166
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/runner/testbench.sv(190) @ 1130: uvm_test_top.env.a.d [DRV] DATA WRITE addr : 10 din : 217
// # KERNEL: UVM_INFO /home/runner/testbench.sv(291) @ 1510: uvm_test_top.env.a.m [MON] DATA WRITE addr:10 data:217
// # KERNEL: UVM_INFO /home/runner/testbench.sv(341) @ 1510: uvm_test_top.env.s [SCO] DATA WRITE OP  addr:10, wdata:217 arr_wr:217
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/runner/testbench.sv(190) @ 1510: uvm_test_top.env.a.d [DRV] DATA WRITE addr : 6 din : 29
// # KERNEL: UVM_INFO /home/runner/testbench.sv(291) @ 1890: uvm_test_top.env.a.m [MON] DATA WRITE addr:6 data:29
// # KERNEL: UVM_INFO /home/runner/testbench.sv(341) @ 1890: uvm_test_top.env.s [SCO] DATA WRITE OP  addr:6, wdata:29 arr_wr:29
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/runner/testbench.sv(190) @ 1890: uvm_test_top.env.a.d [DRV] DATA WRITE addr : 9 din : 125
// # KERNEL: UVM_INFO /home/runner/testbench.sv(291) @ 2270: uvm_test_top.env.a.m [MON] DATA WRITE addr:9 data:125
// # KERNEL: UVM_INFO /home/runner/testbench.sv(341) @ 2270: uvm_test_top.env.s [SCO] DATA WRITE OP  addr:9, wdata:125 arr_wr:125
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/runner/testbench.sv(190) @ 2270: uvm_test_top.env.a.d [DRV] DATA WRITE addr : 3 din : 216
// # KERNEL: UVM_INFO /home/runner/testbench.sv(291) @ 2650: uvm_test_top.env.a.m [MON] DATA WRITE addr:3 data:216
// # KERNEL: UVM_INFO /home/runner/testbench.sv(341) @ 2650: uvm_test_top.env.s [SCO] DATA WRITE OP  addr:3, wdata:216 arr_wr:216
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/runner/testbench.sv(190) @ 2650: uvm_test_top.env.a.d [DRV] DATA WRITE addr : 8 din : 79
// # KERNEL: UVM_INFO /home/runner/testbench.sv(291) @ 3030: uvm_test_top.env.a.m [MON] DATA WRITE addr:8 data:79
// # KERNEL: UVM_INFO /home/runner/testbench.sv(341) @ 3030: uvm_test_top.env.s [SCO] DATA WRITE OP  addr:8, wdata:79 arr_wr:79
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/runner/testbench.sv(190) @ 3030: uvm_test_top.env.a.d [DRV] DATA WRITE addr : 8 din : 215
// # KERNEL: UVM_INFO /home/runner/testbench.sv(291) @ 3410: uvm_test_top.env.a.m [MON] DATA WRITE addr:8 data:215
// # KERNEL: UVM_INFO /home/runner/testbench.sv(341) @ 3410: uvm_test_top.env.s [SCO] DATA WRITE OP  addr:8, wdata:215 arr_wr:215
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/runner/testbench.sv(190) @ 3410: uvm_test_top.env.a.d [DRV] DATA WRITE addr : 1 din : 163
// # KERNEL: UVM_INFO /home/runner/testbench.sv(291) @ 3790: uvm_test_top.env.a.m [MON] DATA WRITE addr:1 data:163
// # KERNEL: UVM_INFO /home/runner/testbench.sv(341) @ 3790: uvm_test_top.env.s [SCO] DATA WRITE OP  addr:1, wdata:163 arr_wr:163
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/runner/testbench.sv(226) @ 4190: uvm_test_top.env.a.d [DRV] DATA READ addr : 2 dout : 0
// # KERNEL: UVM_INFO /home/runner/testbench.sv(311) @ 4190: uvm_test_top.env.a.m [MON] DATA READ addr:2 data:0
// # KERNEL: UVM_INFO /home/runner/testbench.sv(349) @ 4190: uvm_test_top.env.s [SCO] DATA MATCHED : addr:2, rdata:0
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/runner/testbench.sv(226) @ 4590: uvm_test_top.env.a.d [DRV] DATA READ addr : 1 dout : 163
// # KERNEL: UVM_INFO /home/runner/testbench.sv(311) @ 4590: uvm_test_top.env.a.m [MON] DATA READ addr:1 data:163
// # KERNEL: UVM_INFO /home/runner/testbench.sv(349) @ 4590: uvm_test_top.env.s [SCO] DATA MATCHED : addr:1, rdata:163
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/runner/testbench.sv(226) @ 4990: uvm_test_top.env.a.d [DRV] DATA READ addr : 6 dout : 29
// # KERNEL: UVM_INFO /home/runner/testbench.sv(311) @ 4990: uvm_test_top.env.a.m [MON] DATA READ addr:6 data:29
// # KERNEL: UVM_INFO /home/runner/testbench.sv(349) @ 4990: uvm_test_top.env.s [SCO] DATA MATCHED : addr:6, rdata:29
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/runner/testbench.sv(226) @ 5390: uvm_test_top.env.a.d [DRV] DATA READ addr : 7 dout : 0
// # KERNEL: UVM_INFO /home/runner/testbench.sv(311) @ 5390: uvm_test_top.env.a.m [MON] DATA READ addr:7 data:0
// # KERNEL: UVM_INFO /home/runner/testbench.sv(349) @ 5390: uvm_test_top.env.s [SCO] DATA MATCHED : addr:7, rdata:0
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/runner/testbench.sv(226) @ 5790: uvm_test_top.env.a.d [DRV] DATA READ addr : 4 dout : 115
// # KERNEL: UVM_INFO /home/runner/testbench.sv(311) @ 5790: uvm_test_top.env.a.m [MON] DATA READ addr:4 data:115
// # KERNEL: UVM_INFO /home/runner/testbench.sv(349) @ 5790: uvm_test_top.env.s [SCO] DATA MATCHED : addr:4, rdata:115
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/runner/testbench.sv(226) @ 6190: uvm_test_top.env.a.d [DRV] DATA READ addr : 5 dout : 0
// # KERNEL: UVM_INFO /home/runner/testbench.sv(311) @ 6190: uvm_test_top.env.a.m [MON] DATA READ addr:5 data:0
// # KERNEL: UVM_INFO /home/runner/testbench.sv(349) @ 6190: uvm_test_top.env.s [SCO] DATA MATCHED : addr:5, rdata:0
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/runner/testbench.sv(226) @ 6590: uvm_test_top.env.a.d [DRV] DATA READ addr : 3 dout : 216
// # KERNEL: UVM_INFO /home/runner/testbench.sv(311) @ 6590: uvm_test_top.env.a.m [MON] DATA READ addr:3 data:216
// # KERNEL: UVM_INFO /home/runner/testbench.sv(349) @ 6590: uvm_test_top.env.s [SCO] DATA MATCHED : addr:3, rdata:216
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/runner/testbench.sv(226) @ 6990: uvm_test_top.env.a.d [DRV] DATA READ addr : 4 dout : 115
// # KERNEL: UVM_INFO /home/runner/testbench.sv(311) @ 6990: uvm_test_top.env.a.m [MON] DATA READ addr:4 data:115
// # KERNEL: UVM_INFO /home/runner/testbench.sv(349) @ 6990: uvm_test_top.env.s [SCO] DATA MATCHED : addr:4, rdata:115
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/runner/testbench.sv(226) @ 7390: uvm_test_top.env.a.d [DRV] DATA READ addr : 10 dout : 217
// # KERNEL: UVM_INFO /home/runner/testbench.sv(311) @ 7390: uvm_test_top.env.a.m [MON] DATA READ addr:10 data:217
// # KERNEL: UVM_INFO /home/runner/testbench.sv(349) @ 7390: uvm_test_top.env.s [SCO] DATA MATCHED : addr:10, rdata:217
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/runner/testbench.sv(226) @ 7790: uvm_test_top.env.a.d [DRV] DATA READ addr : 7 dout : 0
// # KERNEL: UVM_INFO /home/runner/testbench.sv(311) @ 7790: uvm_test_top.env.a.m [MON] DATA READ addr:7 data:0
// # KERNEL: UVM_INFO /home/runner/testbench.sv(349) @ 7790: uvm_test_top.env.s [SCO] DATA MATCHED : addr:7, rdata:0
// # KERNEL: ----------------------------------------------------------------
// # KERNEL: UVM_INFO /home/build/vlib1/vlib/uvm-1.2/src/base/uvm_objection.svh(1271) @ 7790: reporter [TEST_DONE] 'run' phase is ready to proceed to the 'extract' phase
// # KERNEL: UVM_INFO /home/build/vlib1/vlib/uvm-1.2/src/base/uvm_report_server.svh(869) @ 7790: reporter [UVM/REPORT/SERVER]
// # KERNEL: --- UVM Report Summary ---
// # KERNEL:
// # KERNEL: ** Report counts by severity
// # KERNEL: UVM_INFO :   63
// # KERNEL: UVM_WARNING :    0
// # KERNEL: UVM_ERROR :    0
// # KERNEL: UVM_FATAL :    0
// # KERNEL: ** Report counts by id
// # KERNEL: [DRV]    20
// # KERNEL: [MON]    20
// # KERNEL: [RNTST]     1
// # KERNEL: [SCO]    20
// # KERNEL: [TEST_DONE]     1
// # KERNEL: [UVM/RELNOTES]     1
// # KERNEL:
// # RUNTIME: Info: RUNTIME_0068 uvm_root.svh (521): $finish called.
// # KERNEL: Time: 7790 ns,  Iteration: 62,  Instance: /tb,  Process: @INITIAL#463_2@.
// # KERNEL: stopped at time: 7790 ns
// # VSIM: Simulation has finished. There are no more test vectors to simulate.
// # VSIM: Simulation has finished.
// Done